module cpu(
    // input dos switchs 
    input wire [2:0]op,
    input wire [3:0]D1,
    input wire [3:0]O1,
    in
    
    // input  dos botao key3 e key2
    input botao1,
    input botao2,
    
    // input do lcd
    input EN,
    input RS,
    input WR,
    output reg[7:0] dado,

    input clk,
    output reg[5:0]ledV,
);

parameter loa = ;

always
ope(
op1 = memoria[3]
);


endmodule